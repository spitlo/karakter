module sets

pub const numbers = {
  `A`: '4'
  `B`: '8'
  `C`: ''
  `D`: ''
  `E`: '3'
  `F`: ''
  `G`: '6'
  `H`: ''
  `I`: '1'
  `J`: ''
  `K`: ''
  `L`: ''
  `M`: ''
  `N`: ''
  `O`: '0'
  `P`: ''
  `Q`: ''
  `R`: ''
  `S`: '5'
  `T`: '7'
  `U`: ''
  `V`: ''
  `W`: ''
  `X`: '✕'
  `Y`: ''
  `Z`: '2'
  `a`: '4'
  `b`: '8'
  `c`: ''
  `d`: ''
  `e`: '3'
  `f`: ''
  `g`: '6'
  `h`: ''
  `i`: '1'
  `j`: ''
  `k`: ''
  `l`: ''
  `m`: ''
  `n`: ''
  `o`: '0'
  `p`: ''
  `q`: ''
  `r`: ''
  `s`: '5'
  `t`: '7'
  `u`: ''
  `v`: ''
  `w`: ''
  `x`: '✕'
  `y`: ''
  `z`: '2'
}
