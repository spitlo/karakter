module sets

pub const fairytale = {
  `A`: 'ĄΑЉАдΆ'
  `B`: 'βḂ'
  `C`: 'ĊÇ'
  `D`: 'ĎĐ'
  `E`: 'єξΣЄ'
  `F`: 'Ḟ'
  `G`: 'Ģ'
  `H`: 'њнЂ'
  `I`: 'Ϊ'
  `J`: '⌡'
  `K`: 'ќ'
  `L`: 'ĹĻĽ'
  `M`: 'Ṁ'
  `N`: 'ѝйŅ'
  `O`: 'фθΌ'
  `P`: 'þ'
  `Q`: ''
  `R`: 'Ŕ'
  `S`: 'Ș'
  `T`: '┬†ṪтȚŤ'
  `U`: 'Ů'
  `V`: ''
  `W`: 'Ŵ'
  `X`: 'χЖ'
  `Y`: 'Ų¥Ϋψ'
  `Z`: ''
  `a`: 'ąάαą'
  `b`: 'вБḃ'
  `c`: '¢ς'
  `d`: 'đďδḋ'
  `e`: 'єёē'
  `f`: 'ḟƒ'
  `g`: 'ġ'
  `h`: 'ћђ'
  `i`: 'їΐ'
  `j`: ''
  `k`: ''
  `l`: 'ļľ'
  `m`: 'ṁ'
  `n`: 'ηñņ'
  `o`: 'фоºσ'
  `p`: ''
  `q`: ''
  `r`: 'ѓг'
  `s`: 'ș'
  `t`: 'ṫțł'
  `u`: 'ΰυ'
  `v`: 'ν'
  `w`: 'шώŵ'
  `x`: 'ж'
  `y`: 'џψ'
  `z`: 'ż'
}
