module sets

pub const standard = {
  `A`: 'ĄΑΔΛЉАд▲'
  `B`: '8'
  `C`: '©'
  `D`: 'ĎĐ'
  `E`: 'єξΣΞ3€'
  `F`: ''
  `G`: ''
  `H`: 'њнЂ'
  `I`: 'Ϊ1'
  `J`: ''
  `K`: 'ќк'
  `L`: ''
  `M`: 'м'
  `N`: 'ѝйи'
  `O`: 'фθ0'
  `P`: ''
  `Q`: ''
  `R`: 'яŔ®'
  `S`: 'Ș5'
  `T`: '┬†ṪтȚŤ'
  `U`: ''
  `V`: ''
  `W`: 'Ŵ'
  `X`: 'χ'
  `Y`: 'Ų¥'
  `Z`: ''
  `a`: 'ąάαаą@ª'
  `b`: 'ъьвБ6'
  `c`: '¢'
  `d`: 'đď'
  `e`: 'єё'
  `f`: ''
  `g`: '9'
  `h`: 'ћђ'
  `i`: 'ї'
  `j`: ''
  `k`: ''
  `l`: '1'
  `m`: ''
  `n`: 'η'
  `o`: 'фоº●'
  `p`: ''
  `q`: ''
  `r`: 'ѓг'
  `s`: 'ș'
  `t`: 'ṫțł'
  `u`: ''
  `v`: '▼'
  `w`: 'шώŵ'
  `x`: 'ж×'
  `y`: 'џψ'
  `z`: ''
}
