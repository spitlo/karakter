module sets

pub const cyberpunk = {
  `A`: 'ΔΛА▲4'
  `B`: '8'
  `C`: '©'
  `D`: 'Đ'
  `E`: 'єΣΞ3€'
  `F`: ''
  `G`: ''
  `H`: 'н'
  `I`: '1Ī┃'
  `J`: '⌡'
  `K`: 'к'
  `L`: 'Ľ┕┖'
  `M`: 'м'
  `N`: 'и'
  `O`: 'θ0Ø⓪█'
  `P`: ''
  `Q`: '?'
  `R`: 'Я®'
  `S`: '5$§'
  `T`: '┬†тȚ7'
  `U`: ''
  `V`: '√'
  `W`: 'Ш'
  `X`: 'χ'
  `Y`: 'Ч'
  `Z`: ''
  `a`: 'αа@'
  `b`: 'вБ6'
  `c`: '¢'
  `d`: 'ď'
  `e`: 'є≡'
  `f`: '⌠'
  `g`: '9'
  `h`: 'H'
  `i`: ':īı¡'
  `j`: ''
  `k`: 'κ'
  `l`: '1'
  `m`: ''
  `n`: 'Π∩π'
  `o`: 'о●ø■'
  `p`: ''
  `q`: ''
  `r`: 'гя┍┎'
  `s`: '$'
  `t`: 'Ł┪'
  `u`: 'μ'
  `v`: '▼'
  `w`: 'ш'
  `x`: '×'
  `y`: 'џч'
  `z`: ''
}
