module sets

pub const standard = {
	`A`: 'ĄΑΔΛЉАд▲'
	`B`: '8'
	`C`: '©'
	`D`: 'ĎĐ'
	`E`: 'єξΣΞ3€'
	`F`: ''
	`G`: ''
	`H`: 'њнЂ'
	`I`: 'Ϊ1'
	`J`: ''
	`K`: 'ќк'
	`L`: ''
	`M`: 'м'
	`N`: 'ѝйи'
	`O`: 'фθ0'
	`P`: ''
	`Q`: ''
	`R`: 'яŔ®'
	`S`: 'Ș5'
	`T`: '┬†ṪтȚŤ'
	`U`: ''
	`V`: ''
	`W`: 'Ŵ'
	`X`: 'χ'
	`Y`: 'Ų¥'
	`Z`: ''
	`a`: 'ąάαаą@ª'
	`b`: 'ъьвБ6'
	`c`: '¢'
	`d`: 'đď'
	`e`: 'єё'
	`f`: ''
	`g`: '9'
	`h`: 'ћђ'
	`i`: 'ї'
	`j`: ''
	`k`: ''
	`l`: '1'
	`m`: ''
	`n`: 'η'
	`o`: 'фоº●'
	`p`: ''
	`q`: ''
	`r`: 'ѓг'
	`s`: 'ș'
	`t`: 'ṫțł'
	`u`: ''
	`v`: '▼'
	`w`: 'шώŵ'
	`x`: 'ж×'
	`y`: 'џψ'
	`z`: ''
}

pub const cyberpunk = {
	`A`: 'ΔΛА▲4'
	`B`: '8'
	`C`: '©'
	`D`: 'Đ'
	`E`: 'єΣΞ3€'
	`F`: ''
	`G`: ''
	`H`: 'н'
	`I`: '1Ī┃'
	`J`: '⌡'
	`K`: 'к'
	`L`: 'Ľ┕┖'
	`M`: 'м'
	`N`: 'и'
	`O`: 'θ0Ø⓪█'
	`P`: ''
	`Q`: '?'
	`R`: 'Я®'
	`S`: '5\$§'
	`T`: '┬†тȚ7'
	`U`: ''
	`V`: '√'
	`W`: 'Ш'
	`X`: 'χ'
	`Y`: 'Ч'
	`Z`: ''
	`a`: 'αа@'
	`b`: 'вБ6'
	`c`: '¢'
	`d`: 'ď'
	`e`: 'є≡'
	`f`: '⌠'
	`g`: '9'
	`h`: 'H'
	`i`: ':īı¡'
	`j`: ''
	`k`: 'κ'
	`l`: '1'
	`m`: ''
	`n`: 'Π∩π'
	`o`: 'о●ø■'
	`p`: ''
	`q`: ''
	`r`: 'гя┍┎'
	`s`: '\$'
	`t`: 'Ł┪'
	`u`: 'μ'
	`v`: '▼'
	`w`: 'ш'
	`x`: '×'
	`y`: 'џч'
	`z`: ''
}

pub const fairytale = {
	`A`: 'ĄΑЉАдΆ'
	`B`: 'βḂ'
	`C`: 'ĊÇ'
	`D`: 'ĎĐ'
	`E`: 'єξΣЄ'
	`F`: 'Ḟ'
	`G`: 'Ģ'
	`H`: 'њнЂ'
	`I`: 'Ϊ'
	`J`: '⌡'
	`K`: 'ќ'
	`L`: 'ĹĻĽ'
	`M`: 'Ṁ'
	`N`: 'ѝйŅ'
	`O`: 'фθΌ'
	`P`: 'þ'
	`Q`: ''
	`R`: 'Ŕ'
	`S`: 'Ș'
	`T`: '┬†ṪтȚŤ'
	`U`: 'Ů'
	`V`: ''
	`W`: 'Ŵ'
	`X`: 'χЖ'
	`Y`: 'Ų¥Ϋψ'
	`Z`: ''
	`a`: 'ąάαą'
	`b`: 'вБḃ'
	`c`: '¢ς'
	`d`: 'đďδḋ'
	`e`: 'єёē'
	`f`: 'ḟƒ'
	`g`: 'ġ'
	`h`: 'ћђ'
	`i`: 'їΐ'
	`j`: ''
	`k`: ''
	`l`: 'ļľ'
	`m`: 'ṁ'
	`n`: 'ηñņ'
	`o`: 'фоºσ'
	`p`: ''
	`q`: ''
	`r`: 'ѓг'
	`s`: 'ș'
	`t`: 'ṫțł'
	`u`: 'ΰυ'
	`v`: 'ν'
	`w`: 'шώŵ'
	`x`: 'ж'
	`y`: 'џψ'
	`z`: 'ż'
}
