module sets

pub const loudmouth = {
  `A`: 'Ā'
  `B`: 'β'
  `C`: 'Č'
  `D`: 'Đ'
  `E`: 'Ē'
  `F`: 'Ḟ'
  `G`: ''
  `H`: 'Ħ'
  `I`: 'Ī'
  `J`: ''
  `K`: 'Ќ'
  `L`: ''
  `M`: ''
  `N`: 'П'
  `O`: 'ŌØΘ'
  `P`: 'РṖ'
  `Q`: ''
  `R`: 'Ŕ'
  `S`: 'Ș'
  `T`: 'Ṫ'
  `U`: 'Ū'
  `V`: ''
  `W`: 'Ш'
  `X`: ''
  `Y`: 'Џ'
  `Z`: 'Ż'
  `a`: 'Ā'
  `b`: 'Ḃ'
  `c`: 'Č'
  `d`: 'Đ'
  `e`: 'Ē'
  `f`: 'F'
  `g`: 'G'
  `h`: 'H'
  `i`: 'I'
  `j`: 'J'
  `k`: 'Ќ'
  `l`: 'L'
  `m`: 'M'
  `n`: 'П'
  `o`: 'Ō'
  `p`: 'Р'
  `q`: 'Q'
  `r`: 'Ŕ'
  `s`: 'Ș'
  `t`: 'Ṫ'
  `u`: 'Ū'
  `v`: 'V'
  `w`: 'Ш'
  `x`: 'X'
  `y`: 'Џ'
  `z`: 'Ż'
}
