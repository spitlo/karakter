module sets

pub const moneytalk = {
  `A`: '₳'
  `B`: '฿৳'
  `C`: '₵₡'
  `D`: '₫'
  `E`: '€'
  `F`: '₣'
  `G`: '₲'
  `H`: '₶'
  `I`: '1'
  `J`: 'J'
  `K`: '₭'
  `L`: '£'
  `M`: '₥'
  `N`: '₦₪'
  `O`: '0'
  `P`: '₽₱'
  `Q`: 'Q'
  `R`: '₹'
  `S`: '₷$'
  `T`: '₸₮₺'
  `U`: 'U'
  `V`: 'V'
  `W`: '₩'
  `X`: 'X'
  `Y`: '¥'
  `Z`: '₴'
  `a`: '₳'
  `b`: '฿৳'
  `c`: '₵₡'
  `d`: '₫'
  `e`: '€'
  `f`: '₣'
  `g`: '₲'
  `h`: '₶'
  `i`: '1'
  `j`: 'J'
  `k`: '₭'
  `l`: '£'
  `m`: '₥'
  `n`: '₦₪'
  `o`: '0'
  `p`: '₽₱'
  `q`: 'Q'
  `r`: '₹'
  `s`: '₷$'
  `t`: '₸₮₺'
  `u`: 'U'
  `v`: 'V'
  `w`: '₩'
  `x`: 'X'
  `y`: '¥'
  `z`: '₴'
}
